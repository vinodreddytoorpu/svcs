module simple();
endmodule
